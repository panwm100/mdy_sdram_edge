/*********www.mdy-edu.com ������ƽ� ע�Ϳ�ʼ****************
������רעFPGA��ѵ���о������н�FPGA��Ŀ������Ŀ������Ϳ���������ٷ���̳ѧϰ��http://www.fpgabbs.cn/����������������PCIE��MIPI����Ƶƴ�ӵȼ��������QȺ97925396��������ѧϰ
**********www.mdy-edu.com ������ƽ� ע�ͽ���****************/

module acsii2hex(
    clk     ,
    rst_n   ,
    din     ,
    din_vld ,
    
    dout    ,
    dout_vld    
    );

    parameter      DIN_W =         8;
    parameter      DOUT_W =        4;
    
    input               clk         ;
    input               rst_n       ;
    input [DIN_W-1:0]   din         ;
    input               din_vld     ;

    wire  [DIN_W-1:0]   din         ;
    wire                din_vld     ;

    output[DOUT_W-1:0]  dout        ;
    output              dout_vld    ;

    reg   [DOUT_W-1:0]  dout        ;
    reg                 dout_vld    ;

    always  @(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            dout_vld <= 0;
        end
        else if(din_vld&&((din>=8'd48&&din<8'd58)||(din>=8'd65&&din<8'd71)||(din>=8'd97&&din<8'd103)))begin
            dout_vld <= 1;
        end
        else begin
            dout_vld <= 0;
        end
    end


    always@(posedge clk or negedge rst_n)begin
        if(rst_n==1'b0)begin
            dout <= 0;
        end
        else if(din>=8'd48&&din<8'd58) begin
            dout <= din - 8'd48;
        end
        else if(din>=8'd65&&din<8'd71) begin
            dout <= din - 8'd55;
        end
        else if(din>=8'd97&&din<8'd103) begin
            dout <= din - 8'd87;
        end
        else begin
            dout <= 0;
        end    
    end

    endmodule


